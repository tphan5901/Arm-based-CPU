`include "ALU_Decoder.v"
`include "Main_Decoder.v"

module Control_Unit(Op, RegWrite, ImmSrc, ALUSrc, MemWrite, ResultSrc, Branch, funct3, funct7, ALUControl);

    input[6:0]Op,funct7;
    input[2:0]funct3;
    output RegWrite,ALUSrc,MemWrite,ResultSrc,Branch;
    output[1:0]ImmSrc;
    output[2:0]ALUControl;

    wire[1:0]ALUOp;

    Main_Decoder Main_Decoder(
            .Op(Op),
            .RegWrite(RegWrite),
            .ImmSrc(ImmSrc),
            .MemWrite(MemWrite),
            .ResultSrc(ResultSrc),
            .Branch(Branch),
            .ALUSrc(ALUSrc),
            .ALUOp(ALUOp)
    );
    
    ALU_Decoder ALU_Decoder(

    );


endmodule